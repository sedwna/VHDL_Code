PACKAGE utilities IS
END utilities;

PACKAGE BODY utilities IS

END utilities;